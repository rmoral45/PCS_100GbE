


module one_hot_to_bin
#(
	parameter NB_INPUT  = 20,
	parameter NB_OUTPUT = 
 )