


module block_sync_fsm
#(
 )
 (
 )