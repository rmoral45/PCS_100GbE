`timescale 1ns/100ps

module tb_swap_v2;

localparam NB_DATA = 66;


