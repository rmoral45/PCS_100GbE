module frameGenerator
	#(
	)
	(
		input 
	)